
//`define	CONFIG_SFP_CHECK_OVERFLOW	//溢出检查，适用于正负无穷检查，如果数据永远不超出 ±1.999984741 × ±2^127，则配置为0
//`define	CONFIG_SFP_USE_EXTENDED		//使用扩展精度，接近0的非规约浮点数。不使用为0
