
module convolution
(

);


endmodule


