module conv_core
(
	i_rst,
	i_clk,
	
	i_req,
	i_da,
	
);